// Code your testbench here
// or browse Examples

// `include "mealy_1011_nonoverlap.v"
// `include "mealy_1011_overlap.v"
// `include "moore_1011_nonoverlap.v"
// `include "moore_1011_overlap.v"
// `include "moore_1101_overlap.v"
// `include "mealy_101101_overlap.v"
 `include "mealy_BBCBC_nonoverlap.v"
// `include "moore_BCCB_nonoverlap.v"
// `include "TLController.v"

