//`include "sync_fifo_tb.v"
//`include "async_fifo_tb.v"
`include "async_fifo_grey_tb.v"
//`include "design.sv"


/*PLEASE RUN IN EDA PLAYGROUND (PREFERABLY QUESTASIM SIMULATOR)*/